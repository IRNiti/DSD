-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Tue Dec 01 20:16:07 2015

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY mastermindStatediagram IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        input1 : IN STD_LOGIC := '0';
        input2 : IN STD_LOGIC := '0';
        input3 : IN STD_LOGIC := '0';
        input4 : IN STD_LOGIC := '0';
        output1 : OUT STD_LOGIC
    );
END mastermindStatediagram;

ARCHITECTURE BEHAVIOR OF mastermindStatediagram IS
    TYPE type_fstate IS (state1,state2,state3,state4,state5,state8,state7,state6);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,input1,input2,input3,input4)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state1;
            output1 <= '0';
        ELSE
            output1 <= '0';
            CASE fstate IS
                WHEN state1 =>
                    IF (NOT((input1 = '1'))) THEN
                        reg_fstate <= state1;
                    ELSIF ((input1 = '1')) THEN
                        reg_fstate <= state2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;
                WHEN state2 =>
                    IF ((input2 = '1')) THEN
                        reg_fstate <= state2;
                    ELSIF (NOT((input2 = '1'))) THEN
                        reg_fstate <= state4;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state2;
                    END IF;
                WHEN state3 =>
                    IF ((input2 = '1')) THEN
                        reg_fstate <= state8;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state3;
                    END IF;
                WHEN state4 =>
                    IF ((input3 = '1')) THEN
                        reg_fstate <= state4;
                    ELSIF (NOT((input3 = '1'))) THEN
                        reg_fstate <= state5;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state4;
                    END IF;
                WHEN state5 =>
                    IF (NOT((input3 = '1'))) THEN
                        reg_fstate <= state5;
                    ELSIF ((input3 = '1')) THEN
                        reg_fstate <= state6;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state5;
                    END IF;
                WHEN state8 =>
                    IF (NOT((input2 = '1'))) THEN
                        reg_fstate <= state6;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state8;
                    END IF;

                    IF (NOT((input1 = '1'))) THEN
                        output1 <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        output1 <= '0';
                    END IF;
                WHEN state7 =>
                    IF ((input2 = '1')) THEN
                        reg_fstate <= state3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state7;
                    END IF;
                WHEN state6 =>
                    IF ((input4 = '1')) THEN
                        reg_fstate <= state7;
                    ELSIF (NOT((input4 = '1'))) THEN
                        reg_fstate <= state6;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state6;
                    END IF;
                WHEN OTHERS => 
                    output1 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
